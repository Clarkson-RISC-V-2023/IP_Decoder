module decoder #(
    // Parameters
)(
    // Ports
);

    begin 
        // Logic definition
    end
endmodule;