module tb_decoder #(
    // Parameters
)(
    // No_Ports
);

    begin 
        // Logic definition
    end
endmodule